module onesecond(output reg [0:0] clk, input clk50);
	reg [31:0] counter;
	reg [31:0] delay;
	initial counter = 0;
	initial delay = 25000000;
	initial clk = 1;

	always @(posedge clk50) begin
		counter = counter + 1;
		if (counter > delay) begin
			clk = ~clk;
			counter = 0;
		end
	end
endmodule



//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module ex1(

	//////////// CLOCK //////////
	input 		          		CLOCK2_50,
	input 		          		CLOCK3_50,
	input 		          		CLOCK4_50,
	input 		          		CLOCK_50,

	//////////// SEG7 //////////
	output		 reg    [6:0]		HEX0,
	output		 reg    [6:0]		HEX1,
	output		 reg    [6:0]		HEX2,
	output		 reg    [6:0]		HEX3,
	output		 reg    [6:0]		HEX4,
	output		 reg    [6:0]		HEX5,

	//////////// KEY //////////
	input 		     [3:0]		KEY,

	//////////// SW //////////
	input 		     [9:0]		SW
);

	wire [0:0] sec;
	reg [6:0] digit[9:0]; 
	reg [31:0] t;
	initial t = 0;
	initial begin
		HEX0 = 'h7F;
		HEX1 = 'h7F;
		HEX2 = 'h7F;
		HEX3 = 'h7F;
		HEX4 = 'h7F;
		HEX5 = 'h7F;
		digit[0] = 'h3F; digit[1] = 'h6; digit[2] = 'h5B;
		digit[3] = 'h4F; digit[4] = 'h66; digit[5] = 'h6D;
		digit[6] = 'h7D; digit[7] = 'h7; digit[8] = 'h7F;
		digit[9] = 'h6F;
	end

	onesecond s1(sec, CLOCK_50);

	always @(posedge sec or negedge KEY[0]) begin
		if (!KEY[0])
			t = 0;
		else begin
			if (SW[0])
				t = t+1;
		end
		HEX0 = ~digit[t%10];
		HEX1 = ~digit[(t/10)%6];
		
		HEX3 = ~digit[(t/60)%10];
		HEX4 = ~digit[(t/600)%10];
		HEX5 = ~digit[(t/6000)%10];
	end
endmodule
